                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                  �    (�   ��
   ��:   ���   \U�   \i�   \y�   \y�   jU�   jU�   �_�   \�   ��   ���   ���   ��   �}�  ��V  �uU  �vU  ���  p_�   p}U �\�U �\_ ��p=  � �=  � �  < �         �   ��#   ��*   ���   ���  pU�  pi�  py�  pyU  �UU  �UU  ��   p�   �   �j   �z  ��v  ��u   �u   �u   �u   �w   ��   �?    �5    �=    �?    p5    p5   ��5   ��?   �?                      �    (�   ��
   ��:   ���   \U�   \i�   \y�   \y�   jU�   jU�   �_�   \�   ��   ���   ���  �U=  �yW�  �U��  �U��  ����  �V��  pU��  pU�� �\��? �\�_ ��p=  � �<  � �  < �                                  ?��   �;[U   ���   ���   �W�   ��U   ���U   ?�UU  ���UU  ���U  p��UU  ���UU=   ����  pU��U=  ����U�   ׫~��   �UU��   �VU��   ����   ���_=   ��V}  �p���  �pi��  ���  ��5��  � �   � ��    < �           �:      �:      ���    �VU   �;��    ��_�   k�U�   W�]�   ��]�   �jU�   puUU   p�_U   �uUU   �uU�   ��k�    ��o5    �k�    ����    \U��    \U��    l�u�    ��u=    ���    pUV    �UV     W�      \�      p6      �?     ��?     ��<                            �       ����    ��U�    ���?    ��W�    ;pU�   �;p]�   ��]�   ��_U�   \\U�   _�W�   �?\U�   ��\U�  �W�Z�?   W��_�  \ݯ^U  p���_  �_U�^   lUU�   ����   ����   |���   ��Z�   W_�]   �U��>   �U|?   �� �?   � �   � �   ��?���?��?��<��?��<?���<�<�<�� ��<? <�<�<�<�� ��<� <�?��<��<����<� <��?��<�� ��<� <�<�<��<�� ��? <�<��<��?��?�?��� ��?����?�? � ����?��? � ����?��?0� ��� ?� ?0� ����<<� <��? ����<0�  ��? ����? �  ��? �����? ��?��� ����? ����� ����<0��<���?��<<��<��?�� ?��< �<?���?�?�< �<<���?�?� ���?��?����?� �?�?������ �?�����?��������?����?�?�� ?����?�?��<<����?�?��<0����?��� �? ����?��� ��? ��� ��?��3 �? ����? �3 �<0����? � �<<����? � � ?���� � ��?���?� � ��?��?�?�  � ����?�                                ����������������������������������������������������������������_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_WUUUUUUUUUUUUUUUUUUUUUUUUUUUUե�]UUUUUUUUUUUUUUUUUUUUUUUUUUUUu�_WUUUUUUUUUUUUUUUUUUUUUUUUUUUUե_U����_������WUU��_����W�����U�_U   `5   �5 VUU� X   X   �U�_U   �    6 VUU� �    `   �U�_U   �    6 VUU� �    `   �U�_U   �    6 VUU� �    `   �U�_U   �    6 VUU� �    `����U�_U��� �
 6 VUU� � �� ``UUUU�_U`U��U5 6 VUU� � XU`����U�_U`���U5 6 VUU� � XU�j   �U�_U` ��U5 6 VUU� � XUUU   �U�_U` ��U5 6 VUU� � XUUU   �U�_U` ��U5 6 VUU� � XU�   �U�_U` ��U5 6 VUU� � XU`����U�_U` ` � 6 ���� � �� ``UUUU�_U`��Z    6 6  � �    `����U�_U`UUU    6 6  � �    `   �U�_U`UUU    6 6  � �    `   �U�_U`UUU    6 6  � �    `   �U�_U`UUU5   �5 6  � X   X   �U�_U�jUUU����j�������Z����V�����U�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUU����_��U��W���������_UUUU�_UUUUU   `�U5 � 6  �    XUUUU�_UUUUU   ��U5 6 6  �    XUUUU�_UUUUU   ��U5 6 6  �    XUUUU�_UUUUU   ��U5 6 6  �    XUUUU�_UUUUU����U5 6 ����    XUUUU�_UUUUU`U��U5 6 VUU��
��ZUUUU�_UUUUU����U5 6 ���UU�UUUUUU�_UUUUU   `�U5 6    VU�UUUUUU�_UUUUU   X�U5 6    XU�UUUUUU�_UUUUU   X�U5 6    XU�UUUUUU�_UUUUU   `�U5 �    XU�UUUUUU�_UUUUU����U5 V��� XU�UUUUUU�_UUUUU`U� � VUU� XU�UUUUUU�_UUUUU���    ���� XU�UUUUUU�_UUUUU   �    6  � XU�UUUUUU�_UUUUU   �    6  � XU�UUUUUU�_UUUUU   �    6  � XU�UUUUUU�_UUUUU   `5   �5  � VU�UUUUUU�_UUUUU����Z����j�����UU��UUUUUU�_WUUUUUUUUUUUUUUUUUUUUUUUUUUUUե�]UUUUUUUUUUUUUUUUUUUUUUUUUUUUu�_WUUUUUUUUUUUUUUUUUUUUUUUUUUUUե_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�0��0<<0�3�  �0�3�?�30�                                                                                  �����                              �����                                                               � ��                   �
           �  ��       ?       �         ����� pU5      ��       ��         ����� p�6      pf      �?                    p6�     ���     W�0                  p60     pf     7��                   p6�     ���     7�0                  p�6      pf      ��                    pU5      ��       \5                    ��               �                                                                                                                                                                                                                   �pp�     �
  �  ��  �?  W�  7�  7�  ��  \5  �� ��������� �� �:��?� �
  �  ��  �?  W�  7�  7�  ��  \�  �� _��[��}���� �?       �
  �  ��  �?  W�  7�  7�  ��  _5 ��> ��� ���} ��  �     �
  �  ��  �?  ��  ��  W�  W�  \�  �� _��[��}���� �?       �
  �  ��  �?  ��  ��  W�  W�  \5  �� �V��V��V� �� �:��?� �
  �  ��  �?  ��  ��  W�  W�  _5 ��> �V� �V��W} ��  �     �
  �  ��  �?  _�  W�  W�  [�  l�  �>  {  w  �  �  �:  �?  �*  �? �� ��  |U \ \ l� �V p�  p�  �� �� �� �        �   � ��
 �� �U	 p5 p5 ��
 �[	 �� ��  ��  �� �  �     �
  �  ��  ��  V�  ��  ��  j�  V9  ��  p�  p�  ��  �  �  �  � ��# ��*  �? �U= �p5 �p5 �Z9 ��    � �� ��> �;   ?      �   � ��
 �� `U 0\ 0\ �V `�? ��7  �?  _ �� � �           �
  �  ��  �?  7�  7�  W�  ��  \5 ���������6���>���?        �   ��? ��� ��p�\U��j�^Z?�n�6 ��?[Z��[Z������?��         ��  ��  <<  �/  [�  7�  7�  ��  W�  �>  _� �Z��ii����:��?� ��  ��  <<  �/  [�  7�  7�  ��  W�  ��  _��Z��y���? �?       ��  ��  <<  �/  [�  7�  7�  ��  W�  �> �[� �Z��[m ��  �     ��  ��  �?  �:  ��  ��  W�  W�  W�  �?  _� �Z��ii����:��?� ��  ��  �?  �:  ��  ��  W�  W�  W�  ��  _��Z��y���? �?       ��  ��  �?  �:  ��  ��  W�  W�  W�  �> �[� �Z��[m ��  �     �� �� ��  �� X� W W �U X�  ��  �� pm p] �� ��  ��      �� �� ��  �� X� � W �U X�  �� p� x�5 ��6���;��?     �� �� ��  �� X� � W �U X�  ��  �^ |Z \��������� ���  �3 ��� �Z% ��0 ��0 �U*  W%  � �_ �y �u ��  �  �     ��� ���  �3 ��� �Z% ��0 ��0 �U*  W% �� �^ \Z- ��? ������    ��� ���  �3 ��� �Z% ��0 ��0 �U*  W%  � � �= ��5 ������ ��  �� �<< �/  [�  7� 7�  ��  W� �>  _� �Z��ym����:��?�     �� 0�� �>  �/ 7�0 W�  ��  '� �>0 _� �Z��ym������?� ��  ��  << 
�/�[� 7� (�( ��  W�  �>  �  ��  �� ������� �� ��<<�
�/�[� 7�  �  ��  W�  �>  �  ��  �� ������� ��  ��  <<  �/  [�  ��  ?�  ��  W�  �>  _� �Z��ii����:��?� ��  ��  <<  �/  [�  ��  ?�  ��  W�  ��  _��Z��y���? �?       ��  ��  <<  �/  [�  ��  ?�  ��  W�  �> �[� �Z��[m ��  �     ��  ��  �?  �:  ��  ��  W�  W�  W�  �?  _� �Z��ii����:��?� ��  ��  �?  �:  ��  ��  W�  W�  W�  ��  _��Z��y���? �?       ��  ��  �?  �:  ��  ��  W�  W�  W�  �> �[� �Z��[m ��  �     �� �� ��  �� X� �_ _ �U X�  ��  �� pm p] �� ��  ��      �� �� ��  �� X� �� _ �U X�  �� p� x�5 ��6���;��?     �� �� ��  �� X� �� _ �U X�  ��  �^ |Z \��������� ���  �3 ��� �Z% ��: ��0 �U*  W%  � �_ �y �u ��  �  �     ��� ���  �3 ��� �Z% ��: ��0 �U*  W% �� �^ \Z- ��? ������    ��� ���  �3 ��� �Z% ��: ��0 �U*  W%  � � �= ��5 ������ ��  ��  << ��/ [�  ?�  ?� ��  W�  �> _� �Z��ym����:��?�     �� 0�� �>  �/ ?�0 �  ��  g� �>0 _� �Z��ym������?� ��  ��  << 
�/�[� �� (?�( ��  W�  �>  �  ��  �� ������� �� ��<<�
�/�[� ��  ?�  ��  W�  �>  �  ��  �� ������� ��  ��  <<  �/  \5  <<  |=  �6  p  �>  _� �Z��ii����?�     ��  ��  <<  �/  \5  <<  |=  �6  p=  ��  _��i���? �?           ��  ��  <<  �/  \5  <<  |=  �6  |  �> �W� �_i ��  �         ��  ��  �>  �/  \5  \5  \5  l9  p  �>  _� �Z��ii����?�     ��  ��  �>  �/  \5  \5  \5  l9  p=  ��  _��i���? �?           ��  ��  �>  �/  \5  \5  \5  l9  |  �> �W� �_i ��  �         ��  ��  �?  �:  \9  �5  �5  l=  p  �?  \:  \7  �?  �  �      ��  ��  �?  �:  \9  �5  �5  l=  p  �;  \�  _� ��� ���          ��  ��  �?  �:  \9  �5  �5  l=  `  �>  l�  w� ��� ���          ��  ��  �3  ��  l5  \3  \7  |9  p  �  l5  �5  �  �>  �?      ��  ��  �3  ��  l5  \3  \7  |9  �  �  �5  w�  �� �         ��  ��  �3  ��  l5  \3  \7  |9  p	  �  _9  {�  �� �         ��  ��  <<  �/ �\5 <<  |= �6 �p �>  _� �Z��ii����?�         ��  �� 0�/ �7  << \5� �:  p 0�> _� �Z��ii����?�     ��  ��  << (�/( \5 <<�|=
 �6  p  �>  _� �����������     �� �� << (�/( \5 << |=  �6  p  �>  _� �����������    ������ ?�  �� ����p�p��Z�UU �� �W��^�p~�����:�>�?�?������ ?�  �� ����p�p��Z�UU ���W��^�>p~�?��? �?      ������ ?�  �� ����p�p��Z�UU��� �W��Z��_� ��>  �?    ������ ��  �� �����j�UU�UU�UU �� �W��^�p~�����:�>�?�?������ ��  �� �����j�UU�UU�UU ���W��^�>p~�?��? �?      ������ ��  �� �����j�UU�UU�UU��� �W��Z��_� ��>  �?    ������ ��  ���� �U �U jU VU ��  \� W� W� �� ��  �� ������ ��  ���� �U �U jU VU ��  \� W��W������ 
    ������ ��  ���� �U �U jU VU ��  \� {��y������     ������ �� ��� �V��U� �U� �U� �U�  �� �[5 �z� �v� ���  �:  �� ������ �� ��� �V��U� �U� �U� �U�  �� �[5 �z� �v����� �    ������ �� ��� �V��U� �U� �U� �U�  �� �[5 �V� �^m���� �    ������ ?�  �� ���#�p�pȥZ#�UU�� �W��^�p~�����:�>�?�?    ���̪�3 ?�  �� ����p��UU��j�Ye̫�3�^�p~��{����>�?�?������?����������p#�UU#��Z�UU �� �_�������������>���?���ª��?��
������#�p#�UU��j�UU �� �_�������������>���?                ???333333333333333333????                                ����������������0��������������                                ��������������������������������                                ��������������������������������                                ������������������������������                                �������������������������������                                ������������0���0���0���0���0���                                ��������������������������������                                ��������������������������������                                                                                    ����  �HUU�UU�(P���R�? R� R� R��R�?(P��UU�HUU�H�������    ����,  �lUW�l�^�l5z�l5x�l5x�l5x�l5x�l5x�l�\�lUW�lUUŜ�������    ��<p5����\UU�\��֜��ۜ ۜ ۜ ۜ���\���\UU��o��<p5���    ����  �LUU�L�������0�M90�M90�M90�M90�M9����  �LUU�L�������    ��?�\s5לs9�s9�s9�s9�s9�s9�s9�s9�s9�s9�s9�s9���?�    �����N��l����o�,9��L��L��L��L��L9��<�o��Z�lS�N���������\UU5����'  �'  �'  �'  �'  �'  �'  �'  �'  �'  ؗ���\UU5���              �     ��  h� j��+�������_��[�>��� �� ��        0 �  @�    PU  h� ���+���o����_��[�>��� �� ��                  �  �  �� ����UU����UU����UU��� ��  �?          �  0  �  �  o>  �:  k: �k� ����� �  �                  �  0  �  �  o>  �:  k: �k� ����� �  �� ( �
 
          �  �  �?  �:  ��  ��  ��  �������� ��  
?� ( �      � � 00��<<0k���0K�<d�3d<0I����0l9�?�0���� 3 �           �   ��  γ  r�  �7 0�7 r�  γ  �� �   �                        ���                                    ����                               �����W���                               W�U]�U���                               W�U]�U���                               W�U]�U���                               W�U]�����                               �����W���                               WUUUU����                               �����_���                               WUUUUU���                               WUUUU����           0                   �����_���           0                   WUUUUU���           0                   WUUUU����           0                   �����_���           0                   WUUUUU���           0                   WUUUU����           0                   �����_���           0                   WUUUUU���           0                   WUUUU����           0                   �����_���           �                   WUUUUU���           �                   WUUUU����           �                   �����_���           �                   WUUUUU���           �                  WUUUU����          ��                  �����_���          ��?                  WUUUUU���          ���                  WUUUU����          ���                  �����_���          |��  ����          WUUUUU���          ww�  �UU��          WUUUU����          ww�  �UU��         �����_���         ww�  �����:         WUUUUU���     �� ww�  �ff��:         WUUUU����    �p� ww�  �ff��:         �����_���    �=|= ww�  �ff��:         WUUUUU���    ���� ww�  �ff��:         WUUUU����    p�\� ww�  �ff��:         �����_����   p�\� ww�?  �ff��:         WUUUUU����   �_� ww�?  �ff��:         WUUUU�����   ��_�< ww�?  �ff��?         �����_���� �WU]�3 ww�=  �UU����        WUUUUU����? pU���� ww�=���UU�UUU        WUUUU����߿�pUU]�� ww�=���ffvVUU        �����_���߷������� ww�=���ffv���        WUUUUU���ݿ�pww]�� ww�=���ffv���        WUUUU����ݷ�pww��� ww�=���ffvy]�        �����_���������_�� ww��_��ffvy]�        WUUUUU������pww��� ww�}���gfvy]�   @U  WUUUU����߷�pww]�� ww�}���fvy]�   @D  �����_���߷������� ww�}_��fvy]�   @D  WUUUUU������pww]�� ww�}��?Uuy]�   @D  WUUUU����ݿ�pww���ww�}���sUuy]�   @D  �����_���߷����_��ww�_��sfvy]�   @D  WUUUUU������pww���w�U���fvy]�   @D  WUUUU����ݿ�pww]��w�U���fvy]�   @D  �����_���ݿ�������TwwUw����fvy]�   @D  WUUUUU������pww]��Tw}w?���fvy]�   @D  WUUUU�������|ww������WU�W�fvy]ת��jD  �����_���������3�����_U?sW�gvy]׀���J  WUUUUU����̰w�������w�W�_uy]׀���J  WUUUU��������w�󷶶��_w3W��y]�*���J�����������������|�����_U��W��y]׈����zUUUUUUUUUU������W������w3�UWU}y]ת*����z���������������_U������w��U��}y]ת�����zUUUUUUUUUU����UU���������U��}y]� �����z�������������WUUU���������UWU}y]ת�����zUUUUUUUUUU���_u�U���������U��}��� *����z�������������UUU���������U��}yUU�"����zUUUUUUUUUU������_���������UWU}y�  (�"��������������� \���������U��}y]u�����WuUUUUUUUUUU�����\���������U��}y]u����������������������������������������                                        ����������������������������<��?���������������.�?ο������*⌎ࠈ�������������������������������������������������������������������WUUUUUUUUUUUUU�������    ������?�?�    ����?<<     �� �<<      ��� �<< �    ���<<?�    ����<?     �����<<     ���<��?�    �� <��?�    �WUUUUUUUUUUUUU����������������   0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      0U   0U      ��   ��      ���   ���   �������� �{UUUUU���UUUUU���WUUUUU;����������ծ�����������������,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,�����,��� �,��� �������� 𮪪���� ��������  ���� �             ���   ��   ���   �   ���         �    � ����(      �     �
                                                              �   ��?    ��   �V� ���?�kT����kU�����V���ڿ����Z����:�j����>�UUU���jU�� ����� ����� �����  �����  ����?  ����                         0           �  0           0      �  � 0 ��?   �U�   �� �_T?�kU��������������o�ڿ����Z����:�j����>�UUU���ZUU� ����� ����� �����  �����  ����?  ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���ة������  ��� � � � � �ύ& ��" � t ���d\��]�� � �\����]��� v� ��X�d���# Lq�@H�Z�扭' )��S��� �� �����# �$ �% (z�hX@� ��� Y� ]Ĝ � � � � � � � �* dGdO� ���HdS`�����+� Yĥ$� �%�  ���+�+�&� �������8� ]ĥ1� �2�  ��8�8�3� ¥���J������ Yĥ� �	�  å����� ]ĥ� ��  `����
� _����� |¥S��� a� ��`���ȱ�	ȱ�
ȱ�ȱ�)
��]̅�]̅�)0�ȱ����HȄdd�
� �L¤ ��� �
�� �d��Ȅd���!�"�$ȱ"�%ȱ"�&ȱ"�'ȱ"�()
��]̅)�]̅*�()0�-ȱ"����HȄ!d+d,�&� �� �� �M)��	���d. �`�.�/�1ȱ/�2ȱ/�3ȱ/�4ȱ/�5)
��]̅6�]̅7�5)0�:ȱ/����HȄ.d8d9�3� к� �� �M)��@Ы���d! �������ȱ�ȱ�ȱ�ȱ�)
��]̅�]̅�)0� ȱ����HȄdd�� й� ��� �
�� �d��Ȅd���J
��A̅K�A̅L�K�ȱK�`�J
��G̅K�G̅L�K�ȱK�`H�Z�)?	@�;�;��%;�;����)@��J��;�;��8����)0�Ȅ������d�;� z�h`H�Z�)?	@�;�;��%;�;����)@��J��;�;� �8�� ��)0� Ȅ������d�;� z�h`H�Z�')?	@�;�';��%;�;�,�)��()@��J��;�;�-�8��-��()0�-Ȅ,�)����,�(d,�;� z�h`H�Z�4)?	@�;�4;��%;�;�9�6��5)@��J��;�;�:�8��:��5)0�:Ȅ9�6����9�5d9�;� z�h`� `� `H�Z�H����I���H�O�I)?
���ʅQ��ʅRdP ��z�h`dO�* dG`�P�Q�CȱQ�=ȱQ�>ȱQ�D)
��]̅@�]̅A�D)0�EȄPd?dB�C� ��dS`H�Z�O���LWť=�F�C;�F)��F�B�@��D)@��J��F�F�E�8��E��D)0�EȄB�@����B�DdB�C)�;�I)����
�@����;�;�F�( �;�G��* �G�?�?�>� ��z�h`H�Z�  �   ��dd��� _� |� � `� aĩ��z�h`H�Z�� ��� �dN�M)?�N�D�� �>�N
��M̅"�U̅/�M̅#�U̅0d!d.� ���M)����� ¥M��� �� a�z�h` `�  `�  `�  d� d�8�� �� ��� �� P�� ا      � ��� `�� d�� d��h�� ��h�� ��h�� ا�     ���  2�   ���8��u�����     �\��u��\���� ��� ���\��u��\������8��     � ����� ���8�� �<��     ���h�������     ���������0��1������������0��0�h��     ���0�����h���<�     �|ƚ�|���  �*��x�   �G��G�� �<G�� �G��G�� �G��u-G�� �G��G�� �G���-G��G��8G��G�� �-G��     � �G�� �G�� �<G�� �G�� �G�� �G�� �-G�� �G��G�� �G���-���8G��KG��8G��u-G��8
G��8
G��8
G��K
G��K
G��K
G�� �G��u-G��     � ����� �<�� ����� ���u-�� ����� ����-����8���� �-��     � ��� ��� �<�� ��� ��� ��� �-�� ����� ����-��8��K��8��u-��8
��8
��8
��K
��K
��K
��8��u-��     ��<��D�<���<��D�<���<��D�<��O<��D�<���<��D�<���<��D�<��     �O<��D�<���<��D�<���<��D�<��     ���Ƞ� �  ����   8��� ���� ���� ���� u��� `���     � P��� :��� /��� '��� ��� ���     � �
�� /d��     ���_�����_��     � ��� |�� i�� T�� L�� ?��     �     ����8�S�f�yˀ� 
 O  
 O  
 O  
 O  
 O  
 O  
 O  
 O           / �      �   �  / _      O   �         _         �8   
� �
	 �
�



	�
	

			�
	
	 �
	�

		�
	��tƜ��tƜ��l�~ʜ�B�l����ʇˊ˒ˡ˫�������6̩  � v� �䩁�M �Š b�� ���  � &ک�J [� _Щ  � =� J� �� v� �ש �J [� �� �� �� 
� � .� � [� F� ]ͥ}��������< b�� ����J [� ��L���л��J [� �� b�����L�� v�  ��J [Ţ�(� �Ӣ�(� �ӭ   D� b����L���������i���i���`���}� � �d}L����?�� �����i����0�< b�� ����J [� ��d���}L�͠< b�� ����J [� /Ω�}L�ͥ�������8���إ����}L�ͩ�}` v� �� �ש�t��Z� 0Ϣ	�d� 0ϥ����Z� 0�L΢�c�Z�d��p��s ��抭   D� b�����` v� Q� آ �
�  0Ϣ�\� 0ϩ�c�`�d���i� ��-���n��dy����9ƫ�����y�y�0dy�y��L�����L�Ω 0� b� b� b� b� b�Lf�` v�dt��c��d�	 ���c�(�d�
 ���c�<�d� ���c�P�d� ���c�d�d� ���c�x�d� �楊��(�� 0Ϣ�n�
 0�L&Ϣ�(� 0Ϣ�n�	 0�抭  ���`Zڅ}
e}��qυi�qυp�j�qυs�rdkdl�i
���υXȹ�υY	�)��Y��cz�d m�` (N 		
p�������𮴯��0�p������� v��c�P�d� ���c�\�d� ��d�� b�� ����)���c�P�d� �� b� b�LЩ�c�\�d� �� b� b�   P�	��!���M �ť����� ��d�d�d�d�L��L�̘	�ɿ�˩��M ��慥�)����c�P�d��p��s ��L�� v�dt�ą�����A�G�
��� ��曦������ �� �L{� �� �� b� b� b�  ��� P�ƛ�������� �� �� �� b�  ��L�� P�`�A
mA���х}�c�轞э?轞э@�?�@�} ���A`�A�04�G
mG��Y҅}�c��A�G�YҍE�YҍF�E�F�} ���G` ]!!!!!!!!	5
_    9�AG�GOHI�I�A�B{C�LfNADAEAFAG�V�V�G�H�I(\'\&\%\$\#\"\!\ \\\\\\\\\\\\\\\\\\\\\\
\	\\\\\\\\\ \�\�\�\�\
\	\\\\\\\\\ \�\�\�\�\�\�\c(\'\&\%\$\#\"\!\ \\\\\\\\\\\\\\\\\\\\\\
\	\\\\\\\\\ \�\�\�\�\�\�\�\cZڅ}
e}��:хi�:хp�j�:хs�rdkdl�i
��vхXȹv�	�)��Y���~ep�z���es���~� �� 0��p� 8�~�kdcLe�L���(���cdk��(��(8�~�p��� ��� 0&�$�s� 8倅lddL��ɠ��ddl��Ń�8倅s m�`Zڅ}
e}��:хi�:хp�j�:хs�rdkdl�i
��vхXȹvхY	�)��Y��cz�d m�`H�Z�d�A�ec�T���i �U� � �T��p0���s��z�h` � � 3�`��������(����`�������2��(����`���#�������d��
���������������M ��` �� �� � �� q� b� #�`���"�������d�d�`��)������L��ƥ`���
����� ��`�������� ��d�`�������� ��d�` �� a� 4�`��
��1�T�1�U��jdtddd�d����}�Lե}8��}���}�m�8�}�q���}�L)ե}8��}���}�l�8�}�s��� ��Ti�T�Ui �U���Te��T�Ui �U�d8�x08�(0Ls�dc�m�k�q�pLv�L�եc�(�d8�x08�0L��L�եdes�d��sdlLWթ�8�d�s� �T ��dk�cep�c�(�$0
�(8�c�pL�թ�p�L�եTi�T�Ui �ULv�`H�Z
����X���Y ��z�h`H�ZdX��Y���Z�C�[� � �X�Z��(������%�Zi0�Z�[i �[�Xi(�X�Yi �Y����� ��d�z�h`H�Zd\��]� �\����]�]� ��z�h`d�d�� �t��8��}0�L�֩ 8�}�ndm��qL�֥}�L��8��}�L�֥}�m�8�}�qdn��8��}0�L�֩ 8�}�ddl��sL�֥}�L�֥}8��}�L�֥}�l�8�}�sdd��
e��� �c�(Lץd8�x08�(0L��?L�L�ץn�c�m�k�q�p�c�(�d~�d8�x08� 0��8�d�sLTץdes�d��sdlL�ֽ �}� �ڦ�� ��Lsץ}
�}�~�L`ץ}
�}��  z�dk�~�~�	��cep�c�(�'���pLsש�pLs���L"�`� �c��d�� ��� ��� ���c��d�� ���c��d�� ��#�c��d�� ��`dtdcdddkdl�
����X���Y�(�j�p��s m�`� �c���d�� ��� ��� ���c���d�� ���c���d�� ��#�c���d�� ��`dtdc���ddkdl�
����X���Y�(�j�p��s m�`H�Z
�����X���Y���j ��z�h`H�Z�l� ��Xej�X�Yi �Y���Xek�X�Yi �Y� �Z��[�d� ��Zi(�Z�[i �[���Zec�Z�[i �[� � ڱX�t� ���1Z�
��Z�QZ�Z��p�����s��Zi(�Z�[i �[�Xej�X�Yi �Y��z�h`��t��j� �
��W�TȹW�Udkdl��p��s���L�8�
��T�XȱT�Y���~i�����i����i(����i����~Ś��Ś08嚅p���8�~�kdcL��L�ń��8嚅cdk�ń0��8�~�p8��L�٩�p��ś���ś088囅s�1��8倅lddL�Ņ�!8囅ddl��Ń�8倅s8��Lک�s ����
�dt��L>�`d�d�d�d�d�dߩ ������`� ������d�`dudvdwdzdyd{d|���d�d�d�d�����P����
��5�T�5�U� � �T� �Ti�T�Ui �U��?�L}ڥ�

�� ��癜 ������ � �虧 �虲 �����d�d�d���

��'腭�'腸�'腮�'腹`dudvdwdzdyd{d|d���d�d�d�d��������P����

�� ��癜 ������ � �虧 �虲 �����d�d�d�d�d�d�d�d�d�d���

��'腭�'腸�'腮�'腹����`H�Z�l� ��Xej�X�Yi �Y���Xek�X�Yi �Y� �Z�@�[�d� ��Zi0�Z�[i �[���Zec�Z�[i �[� � ڱX�t� ���1Z�
��Z�QZ�Z��p�����s��Zi0�Z�[i �[�Xej�X�Yi �Y��z�h`����d}d�L#�8��}�}J��春���d}d�L>�8��}�}JJJ��早 �}���
�}i�}�������Lp�8����}�}Lp�8����}��~���	8�~j�~����}� �%~� ��
��M �� �� ��`���ei�f���gi�h �� 2�  �`���@���~i�����i�� �ݥ}�'d�d�d���冦�
�񥭅������'�} ީ��M ��`���-���~i�����i�� �ݥ}�d�d穀�M �����i���`� ���$� ���~i�����i�� �ݥ}� ����������`���L�ݥ��ei�f���gi�h� ���+���%���~i�����i�� �ݥ}���������(������`H�Z�e�~���
�"�f�~���gŀ�Ń�
��hŀ�����}�� �}� z�h`�����i �ݥ�i �ޥ�i ���`���e}�ޥ�i ���`�u��u�v��v�w��w�  ������L����- D� ����c��d� �� b� b�   D����� �J [�L����L�̊	����C��i�����} =�}���, ���z�z�0dz�zi����i(8��暥��0���L�ߊ	����>��8������} =�}���� ���y�y�0dy�yi
����8��

ƚ��� d�L�ߊ	����A��8������} �}���* ���{�{�0d{�{i����8����8���� d�L�ߊ	����A��i�����} �}���- ���|�|�0d|�|i����i_8���i���D0�D���	���� �ृ���uL�ߊ	���� �ृ���v`��)��	�����L��ƫL���
8�����L����i��`��)��	����
��8���L���i��L���ƫL��`��JJJJ�~��JJ���)���L9����L9� �}L<� g�`��JJ���JJJJ�~��)�0�0�~Lc� �}Lf� g�`ڥ�
��1�T�1�U�~��Ti�T�Ui �U���Te�T�Ui �U� �T� �� �}�`d�������������������������`d����!����8�����ة
����������������`����������d�d�`�����L�Ƣ`������
����d�d�`� �������	����� ��`��������LG�֜����`H�Z��)�L�᥂JJJJ�~�nJJ��n)�� �}Lw� ��z�h`H�Z��)�L�᥁JJ��oJJJJ�~�o)�� �}L�� ��z�h`H�Z��
��1�T�1�U�~��Ti�T�Ui �U���Te�T�Ui �U� �T� �� �}L�� ��z�h`H���5���ei�f���gi�h���~i�����i�� �ݥ}�� �}����}h`� ���8��ɵ��LI���LI�d�d�d�d�d����n���o���Ƅ愵�e�)� �!�o8����n�����} M�}��������L����!�ni���o�����} {�}���P�����L����!�oi���n�����} M�}���+�����L�����n8����o�����} {�}�������效� �L_⥕�L��i)�� R�LI䥕��%���� L:㥔��L:㥒��L:��� R�LI���C���报�)�� ��L�㥔�报�)����L�㥒�报�)����L���� R�LI� �ɥnū[�oŶ.���#���
��� R�LI�报�)�L���� R�LI䥒��LF㥔����L��报�)�L�� �� R�LI䥑��LF�oŶ.���#���
��� R�LI�报�)�L���� R�LI䥒��LF㥓����L��报�)�L�� �� R�LI䥑��LF����L0�`H�Z� ���i��� ��i����8���L������i��� ��i
����i��L������i��� ��i����i��L������i��� ��i����8���z�h`H�Z����� ����b��a� �e���g�g�d�e�c ��g�r� ��g��d�f���h�g�g�d�e�c� ����a ���h�h�h�d�f�c��a��� ��h�D� �L� � �g�d��a�e�c� �� ��ei�e�c ��f�c��� ��f8��f�c ��f�T� �LW�z�h`xH�Z��
���\��	�)��]�a�}�b�~�d�A�^���_�cJJ��\%��^�\i�\�]i �]�~�~� �Ȁ��}�}� ��b�~�L��z�hX`H� �� �����h`H�Z�/���� ���� ��z�h` @�@H�Z




���)�& z�h`H�  ���� P�h`Hڭ  �����h`Hd��  ������0�h`�Z�P���� ���� ��z�`H�Zd\�@�]� � � �\����]���z�h`H�Z
���煆载煇� ���$��a��b��c��d�8�7�` ��Ȁ�z�h`H�Z�)�JJJJ�` ��)�` ��z�h`xH�Z�`�a��$��b��%��c��&��d��'�����\����]��}�d�A�^���_�c�\�^�\Ȳ\�^�\��}���c�cz�hX`aaTOP$SCORE$STAGE$ada$GAMEaOVER$PAUSE$START$CONTINUE$END$PROGRAMEaBY$aaLIHONG$aGRAPHaaaBY$aaZHANGLIa$aMUSICaaaBY$aXIAOLIWEI$A�G�M�S�W�a�g�m�v�z������p����0�p���𜠅��        ,�,�PP0� `�p$pP$�0pp$P(P�P00�0p0�m���������!�!�#���0�p�����0�p�����0�p�����0�p�����0�p�����0�p�����0�p�����0�p����0�p����0�p����0�p����0�p����0�p����0�p����0�p����0�p����0�p����0�p����0�����0�p�����0�p�����0�p�����0�p�����0�  0@P`p��I����D����?����:����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         M����
�I�����E�������������������������������������������������������������� �� �� �� �� �� �� �� �� �� �� ����������������������������� � � ���������������� � � �������������������������������������������������8 � ������������������������������������������������������ ��8���������  �  �  �����  �  �  ���  �  �  �����  �  �  ���  �  �  ��������������������� ��8���������� �� �� ���������������������������  �  �  �������������������?�������������������������� �� �� �� �� �� �� ������������������������������������������� �  �  � ���� � � ��� �  �  � �����������������  �  �  �����  �  �  ���  �  �  �����  �  �  ���  �  �  ��������� �� �� ��� �� �� ����� �� �� ����� �� �� ����� �� �� ��� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P�� 0`��� P�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____^^^^^^____^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             T� �U�